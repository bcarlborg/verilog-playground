`ifndef DECODER_4TO16_V
`define DECODER_4TO16_V

module decoder_4to16(
  input [3:0] in,
  output [15:0] out
);

  assign out = in[3] & in[2] & in[1] & in[0] ? 16'b1000000000000000
            : in[3] & in[2] & in[1] & ~in[0] ? 16'b0100000000000000
            : in[3] & in[2] & ~in[1] & in[0] ? 16'b0010000000000000
            : in[3] & in[2] & ~in[1] & ~in[0] ? 16'b0001000000000000
            : in[3] & ~in[2] & in[1] & in[0] ? 16'b0000100000000000
            : in[3] & ~in[2] & in[1] & ~in[0] ? 16'b0000010000000000
            : in[3] & ~in[2] & ~in[1] & in[0] ? 16'b0000001000000000
            : in[3] & ~in[2] & ~in[1] & ~in[0] ? 16'b0000000100000000
            : in[2] & in[1] & in[0] ? 16'b0000000010000000
            : in[2] & in[1] & ~in[0] ? 16'b0000000001000000
            : in[2] & ~in[1] & in[0] ? 16'b0000000000100000
            : in[2] & ~in[1] & ~in[0] ? 16'b0000000000010000
            : in[1] & in[0] ? 16'b0000000000001000
            : in[1] & ~in[0] ? 16'b0000000000000100
            : in[0] ? 16'b0000000000000010
            : 16'b0000000000000001;
endmodule

`endif
